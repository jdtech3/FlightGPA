module FlightGPA ();

endmodule